module alu4 (
    input                       clk,
    input                       rst,

    input           [2: 0]      sel,
    input           [3: 0]      A,
    input           [3: 0]      B,
    output reg      [3: 0]      C
);
    
endmodule