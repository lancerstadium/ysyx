    module convLayerMultiTB();
    parameter   DATA_WIDTH              = 16;                   // Data width
    parameter   FLOAT_MODE              = 1;                    // 0: SInt, 1: Float
    parameter   D                       = 1;                    // fit depth
    parameter   S                       = 5;                    // fit size
    parameter   H                       = 32;                   // img height
    parameter   W                       = 32;                   // img width
    parameter   K                       = 6;                    // Number of fits applied
    reg                                 clk, rst;               // Signal
    reg         [D*H*W*DATA_WIDTH-1: 0] img;                    // We test with a 1*32*32 img
    reg         [K*D*S*S*DATA_WIDTH-1: 0] fits;                 // 6 fits with dimensions: Depth:1 Height:5 and Width:5
    wire        [K*(H-S+1)*(W-S+1)*DATA_WIDTH-1:0] res;

    localparam PERIOD = 100;

    integer i, rCnt;

    always
        #(PERIOD/2) clk = ~clk;
        
        
    initial begin 
        #0
        clk = 1'b0;
        rst = 1;
        //We test with a padded img and the filter of the first convolution layers
        img = 16384'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000326638fd3bf038fd32460000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000032063b773be83be83be83b6f000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000032c73b1f3bf03be83b7f3b4f3be833272606000000000000000000000000000000000000000000000000000000000000000000000000000000000000290533883b073be83bf03be83a5635453be83bf037a8000000000000000000000000000000000000000000000000000000000000000000000000000000000000391d3be83be83be83bf03be83be8360639ee3bf0393d0000000000000000000000000000000000000000000000000000000000000000000000000000000032663b773bf03bf039f637273bf03b2731e634f53c003945000000000000000000000000000000000000000000000000000000000000000000000000000032063b773be83be8399e2a0634b537982d45000000003bf03ba032460000000000000000000000000000000000000000000000000000000000000000000030c5392d3bf03b4f3a8735450000000000000000000000003bf03be8392d0000000000000000000000000000000000000000000000000000000000000000270739963be83b8834742cc52f070000000000000000000000003bf03be83a1e000000000000000000000000000000000000000000000000000000000000000033273be83be833e80000000000000000000000000000000000003bf03be83a1e00000000000000000000000000000000000000000000000000000000000000003a363bf039f600000000000000000000000000000000000000003c003bf03a2600000000000000000000000000000000000000000000000000000000000034c53bb83be8370700000000000000000000000000000000000000003bf03be838a500000000000000000000000000000000000000000000000000000000000035553be83b372e46000000000000000000000000000000002707383c3bf039d62a0600000000000000000000000000000000000000000000000000000000000035553be83aff000000000000000000000000000000002707381c3be83b0f3474000000000000000000000000000000000000000000000000000000000000000035553be8388d00000000000000000000000000003206392d3be8396d00000000000000000000000000000000000000000000000000000000000000000000000035653bf03b0f00000000000000000000000037273b773bf03915000000000000000000000000000000000000000000000000000000000000000000000000000035553be83bd0389532062f47355539963b0f3bf03aff393d3307000000000000000000000000000000000000000000000000000000000000000000000000000035553be83be83be83b2f3abf3be83be83be83a2638140000000000000000000000000000000000000000000000000000000000000000000000000000000000002f073a3e3be83be83bf03be83be83b4f388d0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002e4638043be83bf03be8386c30a50000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        fits[0*S*S*DATA_WIDTH+:S*S*DATA_WIDTH] = 400'h346b33f83146351432de310e2cc624deb409b3a2b61ab4c8b679b63bb455b48d2b45b08b2bdbb4c0b536b4b9b598b810b521;
        fits[1*S*S*DATA_WIDTH+:S*S*DATA_WIDTH] = 400'h2beb2d7b319a3303349830989e6132afa8af343b345632da34043406345c30ebac9dacf7b0ec2464b26d2e3bb2c4b33cb203;
        fits[2*S*S*DATA_WIDTH+:S*S*DATA_WIDTH] = 400'ha610312fad4522feac2330d832a4319ba5ecaac229349a10afb12f4aaeb8aadb2f99b26021bdac24a968aef7321c29c82d35;
        fits[3*S*S*DATA_WIDTH+:S*S*DATA_WIDTH] = 400'h240634542fc9375033bf3851365635c4a3bd2b162aac2a602c7e31812d6a35d03782310c37c130e932e22624a6b8ab7da1f3;
        fits[4*S*S*DATA_WIDTH+:S*S*DATA_WIDTH] = 400'ha99baabc2aa33113af6bb1db23c8aa0ab69ab575b6ebb60e16d4b1dfac5a31be2f9c2b2ab298b1b6b2cdae2db5c6b4f0af69;
        fits[5*S*S*DATA_WIDTH+:S*S*DATA_WIDTH] = 400'h37fe37f0380b340434572f01309f31f32e76a6dd2aba9fa734cf303536562c91338e34322f47b1442217a6c2a8eba2a8addc;
        $display("[img]: ");
        for (i = H*W-1; i >=0; i = i - 1) begin
            $write(" %h", img[i*DATA_WIDTH+:DATA_WIDTH]);
            if(i % (W) == 0)begin
                $display(""); 
            end
        end
        rCnt = 0;
        $display("[fit%2d]: ", rCnt);
        for (i = K*S*S-1; i >=0; i = i - 1) begin
            $write(" %h", fits[i*DATA_WIDTH+:DATA_WIDTH]);
            if(i % (S) == 0) begin
                $display("");
                if(i % (S*S) == 0 && i != 0) begin
                    rCnt = rCnt + 1;
                    $display("[fit%2d]: ", rCnt);
                end
            end
        end
        #(PERIOD)

        rst = 0;
        
        #(7*1457*PERIOD)  // we wait for extra clock cycles to prove that the result does not change with extra clock cycles can be used in pipelining
        rCnt = 0;
        $display("[res%2d]: ", rCnt);
        for (i = K*(H-S+1)*(W-S+1)-1; i >=0; i = i - 1) begin
            $write(" %h", res[i*DATA_WIDTH+:DATA_WIDTH]);
            if(i % (W-S+1) == 0) begin
                $display("");
                if(i % ((H-S+1)*(W-S+1)) == 0 && i != 0) begin
                    rCnt = rCnt + 1;
                    $display("[res%2d]: ", rCnt);
                end
            end
        end
        $finish;
    end

    convLayerMulti#(
        .DATA_WIDTH(DATA_WIDTH),
        .FLOAT_MODE(FLOAT_MODE),
        .D(D),
        .S(S),
        .H(H),
        .W(W),
        .K(K)
    ) UUT (
        .clk(clk),
        .rst(rst),
        .img(img),
        .fits(fits),
        .res(res)
    );

endmodule
