module tanh #(
    parameter   DATA_WIDTH              = 32                    // Data width, default: 32 bits
) (
    input       [DATA_WIDTH - 1: 0]     X,                      // F16/32/64: X
    output reg  [DATA_WIDTH - 1: 0]     Y                       // F16/32/64: Y
);



endmodule