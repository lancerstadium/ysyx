module procElemTB();

    reg clk, rst;
    reg [31:0] A, B, R;
    wire [31:0] C;

    localparam PERIOD = 100;

    always
        #(PERIOD/2) clk = ~clk;

    // A = 11000010101111011011110100010100, B = 11000011000010001100111111100110, C = 01000110010010101100110100010001
    // A =    -94.869, B =   -136.812, C =    12979.268, C_hw =    12979.267, Bias =    0.001
    // A = 11000010111101110101101000010000, B = 11000010110000011101010111000111, C = 01000110110000110000101101000010
    // A =   -123.676, B =    -96.918, C =    24965.631, C_hw =    24965.629, Bias =    0.002
    // A = 01000001010001000110110111110000, B = 01000011000000000001101100111000, C = 01000110110011110101010010111101
    // A =     12.277, B =    128.106, C =    26538.371, C_hw =    26538.369, Bias =    0.002
    // A = 01000001110001001111001010010000, B = 11000011001100010101010001010100, C = 01000110101011010011100110011000
    // A =     24.618, B =   -177.329, C =    22172.797, C_hw =    22172.797, Bias =    0.000
    // A = 01000010111011010001100011011000, B = 11000011000100111110001010110110, C = 01000101100100010000100101110000
    // A =    118.549, B =   -147.886, C =     4641.178, C_hw =     4641.180, Bias =   -0.002
    // A = 11000011001101111111011111111000, B = 01000010100001000001001001111000, C = 11000101111010101001101100010110
    // A =   -183.969, B =     66.036, C =    -7507.388, C_hw =    -7507.386, Bias =   -0.002
    // A = 01000010001100111011001100011000, B = 11000010000001000110101110001000, C = 11000110000011001000101001111111
    // A =     44.925, B =    -33.105, C =    -8994.627, C_hw =    -8994.624, Bias =   -0.003
    // A = 01000011001100011001000101110000, B = 01000011000000100101100011010110, C = 01000110010111010001101101100110
    // A =    177.568, B =    130.347, C =    14150.848, C_hw =    14150.850, Bias =   -0.002
    // A = 11000010011010100011011101011000, B = 01000010101000010110000110001000, C = 01000110000100110100100001100010
    // A =    -58.554, B =     80.690, C =     9426.093, C_hw =     9426.096, Bias =   -0.003
    // A = 11000010111101011110111010110011, B = 11000001110000011000011000010000, C = 01000110010000011100001011010001
    // A =   -122.966, B =    -24.190, C =    12400.702, C_hw =    12400.704, Bias =   -0.002
    // A = 01000010100111110011111110011100, B = 01000010101101111111110011011100, C = 01000110100110100001101101001010
    // A =     79.624, B =     91.994, C =    19725.645, C_hw =    19725.645, Bias =    0.000
    // A = 01000010101100101001010110000100, B = 11000011001001111100100101101100, C = 01000101100101000011110011111100
    // A =     89.292, B =   -167.787, C =     4743.621, C_hw =     4743.623, Bias =   -0.002
    // A = 11000010100111101111111010010101, B = 11000010010011110000011101000100, C = 01000110000010100110100010101100
    // A =    -79.497, B =    -51.757, C =     8858.167, C_hw =     8858.168, Bias =   -0.001
    // A = 01000011000110001010001000011000, B = 11000000110000111010011110000000, C = 01000101111101111010011110000100
    // A =    152.633, B =     -6.114, C =     7924.938, C_hw =     7924.939, Bias =   -0.002
    // A = 01000010010001111100100101110100, B = 11000010110110111111000101111101, C = 01000101000110000000001101110000
    // A =     49.947, B =   -109.972, C =     2432.213, C_hw =     2432.215, Bias =   -0.002
    // A = 00111110100000110000001000000000, B = 01000011000110110001001111010010, C = 01000101000110100111111001010010
    // A =      0.256, B =    155.077, C =     2471.893, C_hw =     2471.895, Bias =   -0.002
    // A = 11000010001110110010001010010000, B = 01000010100110010010100011110100, C = 11000100100010101101100110111010
    // A =    -46.784, B =     76.580, C =    -1110.806, C_hw =    -1110.804, Bias =   -0.002
    // A = 11000011000011011101011100010000, B = 01000011001001010111111000111010, C = 11000110110000000001000010110101
    // A =   -141.840, B =    165.493, C =   -24584.359, C_hw =   -24584.354, Bias =   -0.006
    // A = 01000000100101011111011001000000, B = 01000010101001011000111010000100, C = 11000110101111010000100011011100
    // A =      4.686, B =     82.778, C =   -24196.434, C_hw =   -24196.430, Bias =   -0.004
    // A = 01000011001111000010100111101000, B = 11000010100110011000011111000110, C = 11000111000101101111000011011001
    // A =    188.164, B =    -76.765, C =   -38640.855, C_hw =   -38640.848, Bias =   -0.008

    initial begin
        #0
        clk = 1'b0;
        rst = 1;
        // A = 2 , B = 3
        A = 32'b11000010101111011011110100010100;
        B = 32'b11000011000010001100111111100110;
        R = 32'b01000110010010101100110100010001;

        #(PERIOD/4)
        rst = 0;

        #(PERIOD/2)
        $display("A = %b, B = %b, C = %b, Bias = %b", A, B, C, C ^ R);

        // A = 1 , B = 5
        #(3*PERIOD/4)
        A = 32'b01000001010001000110110111110000;
        B = 32'b01000011000000000001101100111000;
        R = 32'b01000110110011110101010010111101;

        #(4*PERIOD/5)
        $display("A = %b, B = %b, C = %b, Bias = %b", A, B, C, C ^ R);

        #(PERIOD)
        $finish;
    end

    procElem PE (
        .clk(clk),
        .rst(rst),
        .A(A),
        .B(B),
        .C(C)
    );

endmodule
